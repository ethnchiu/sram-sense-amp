** sch_path: /foss/designs/sram-sense-amp/xschem/sram-sense-amp.sch
**.subckt sram-sense-amp
V1 VDD GND {VDD}
V2 BLB GND {VDD - dv}
V3 BL GND {VDD}
V4 SE GND PULSE(0 {VDD} 2n 10p 10p 2n 5n)
XM8 net3 SE GND GND sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM9 OUT net2 VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM1 net1 BLB net3 GND sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM4 net3 BL net2 GND sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM3 net2 net1 VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM2 VDD net1 net1 VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM6 OUT net2 GND GND sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
**** begin user architecture code


.lib cornerMOSlv.lib mos_tt

.param VDD=1.2
.param dv=0.02

.tran 0.1p 10n

.control
run
set wr_singlescale
set wr_vecnames
wrdata data.txt v(BL) v(BLB) v(SE) v(OUT)
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
